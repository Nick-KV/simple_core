library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package test_pkg is

	constant r_file1_c : string := "../../../../../sim/mif/inp1_tb.mif";
	constant r_file2_c : string := "../../../../../sim/mif/inp2_tb.mif";
	constant r_file3_c : string := "../../../../../sim/mif/inp3_tb.mif";
	constant r_file4_c : string := "../../../../../sim/mif/inp4_tb.mif";
	constant r_file5_c : string := "../../../../../sim/mif/inp5_tb.mif";
	constant w_file1_c : string := "../../../../../sim/mif/out1_tb.mif";
	constant w_file2_c : string := "../../../../../sim/mif/out2_tb.mif";
	constant w_file3_c : string := "../../../../../sim/mif/out3_tb.mif";
	constant w_file4_c : string := "../../../../../sim/mif/out4_tb.mif";
	constant w_file5_c : string := "../../../../../sim/mif/out5_tb.mif";
	
end test_pkg;

package body test_pkg is

end test_pkg;